module cpu (...); // simplified top-level CPU module endmodule
