module pipelined_cpu (
    input clk,
    input reset
);
// Just a placeholder — will connect IF → ID → EX → MEM → WB stages in future
endmodule
